module test(
    input a,
    output b // adding "reg"
);
    assign b=a;
endmodule