`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/11/08 21:09:41
// Design Name: 
// Module Name: testbench_source_q5
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module testbench_source_q4();
    reg [2:0] x;
    reg [2:0] e;
    wire [7:0] y;

	
    mux mux_test(x,e,y);
	
    initial begin
            x = 3'b000; e = 3'b000;
            #10	x = 3'b001; e = 3'b000;
			#10	x = 3'b010; e = 3'b000;
			#10	x = 3'b011; e = 3'b000;
			#10	x = 3'b100; e = 3'b000;
			#10	x = 3'b101; e = 3'b000;
			#10	x = 3'b110; e = 3'b000;
            #10	x = 3'b111; e = 3'b000;

            #10	x = 3'b000; e = 3'b001;
            #10	x = 3'b001; e = 3'b001;
			#10	x = 3'b010; e = 3'b001;
			#10	x = 3'b011; e = 3'b001;
			#10	x = 3'b100; e = 3'b001;
			#10	x = 3'b101; e = 3'b001;
			#10	x = 3'b110; e = 3'b001;
            #10	x = 3'b111; e = 3'b001;
            
            #10	x = 3'b000; e = 3'b010;
            #10	x = 3'b001; e = 3'b010;
			#10	x = 3'b010; e = 3'b010;
			#10	x = 3'b011; e = 3'b010;
			#10	x = 3'b100; e = 3'b010;
			#10	x = 3'b101; e = 3'b010;
			#10	x = 3'b110; e = 3'b010;
            #10	x = 3'b111; e = 3'b010;
            
            #10	x = 3'b000; e = 3'b011;
            #10	x = 3'b001; e = 3'b011;
			#10	x = 3'b010; e = 3'b011;
			#10	x = 3'b011; e = 3'b011;
			#10	x = 3'b100; e = 3'b011;
			#10	x = 3'b101; e = 3'b011;
			#10	x = 3'b110; e = 3'b011;
            #10	x = 3'b111; e = 3'b011;
            
            #10	x = 3'b000; e = 3'b100;
            #10	x = 3'b001; e = 3'b100;
			#10	x = 3'b010; e = 3'b100;
			#10	x = 3'b011; e = 3'b100;
			#10	x = 3'b100; e = 3'b100;
			#10	x = 3'b101; e = 3'b100;
			#10	x = 3'b110; e = 3'b100;
            #10	x = 3'b111; e = 3'b100;

            #10	x = 3'b000; e = 3'b101;
            #10	x = 3'b001; e = 3'b101;
			#10	x = 3'b010; e = 3'b101;
			#10	x = 3'b011; e = 3'b101;
			#10	x = 3'b100; e = 3'b101;
			#10	x = 3'b101; e = 3'b101;
			#10	x = 3'b110; e = 3'b101;
            #10	x = 3'b111; e = 3'b101;

            #10	x = 3'b000; e = 3'b110;
            #10	x = 3'b001; e = 3'b110;
			#10	x = 3'b010; e = 3'b110;
			#10	x = 3'b011; e = 3'b110;
			#10	x = 3'b100; e = 3'b110;
			#10	x = 3'b101; e = 3'b110;
			#10	x = 3'b110; e = 3'b110;
            #10	x = 3'b111; e = 3'b110;

            #10	x = 3'b000; e = 3'b111;
            #10	x = 3'b001; e = 3'b111;
			#10	x = 3'b010; e = 3'b111;
			#10	x = 3'b011; e = 3'b111;
			#10	x = 3'b100; e = 3'b111;
			#10	x = 3'b101; e = 3'b111;
			#10	x = 3'b110; e = 3'b111;
            #10	x = 3'b111; e = 3'b111;

    end
endmodule
